module ifetch(
	input logic clk, reset, StallF,
	input logic [31:0] PC,	// Next PC value
	output logic [31:0] PCF, PCPlus4F);

//	flopr #(32) IFReg(clk, reset, PC, PCF);
        always_ff @(posedge clk, posedge reset)
          if (StallF);
          else if (reset) PCF <= 32'b0;
          else PCF <= PC;
	adder #(32) IFAdd(PCF, 32'b100, PCPlus4F);

endmodule
