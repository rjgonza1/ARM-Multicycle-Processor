dlfkajds;flsdj
